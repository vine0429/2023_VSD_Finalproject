`define CPU_CYCLE     7.0 // 100Mhz
`define MAX           3000000 // 3000000
