`define CPU_CYCLE     5.8 // 100Mhz
`define MAX           3000000 // 3000000
