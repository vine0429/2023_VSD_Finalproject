`define CPU_CYCLE     7.0 // 100Mhz
`define MAX           6000000 // 3000000
`define AXI_CYCLE     25.0 // 40Mhz
