`define CPU_CYCLE     6.0 // 100Mhz
`define MAX           30000000 // 3000000
`define AXI_CYCLE     25.0 // 40Mhz
