
`define FRAME_WIDTH  640 
`define FRAME_HEIGHT 320
`define ROW_MB_NUM FRAME_WIDTH >> 4
`define FRAME_WIDTH_DIV4  FRAME_WIDTH >> 2
`define FRAME_HEIGHT_DIV4 FRAME_HEIGHT >> 2
